// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_UUT_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_UUT_AXI_ID_W 4
`define IOB_UUT_AXI_LEN_W 8
`define IOB_UUT_AXI_ADDR_W 18
`define IOB_UUT_AXI_DATA_W 32
`define IOB_UUT_BAUD 3000000
`define IOB_UUT_FREQ 100000000
`define IOB_UUT_SIMULATION 1
