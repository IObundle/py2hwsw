// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_AXI_ID_W 4
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_AXI_LEN_W 8
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_AXI_ADDR_W 30
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_AXI_DATA_W 32
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_BAUD 115200
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_FREQ 100000000
`define IOB_UART_TESTER_IOB_AES_KU040_DB_G_XILINX 1
