// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_dma_csrs.vh"
`include "iob_dma_csrs_conf.vh"
`define IOB_CSRS_ADDR_W `IOB_DMA_CSRS_ADDR_W
