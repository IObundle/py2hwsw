// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UART_DATA_W 32
// Core Configuration Macros.
`define IOB_UART_RST_POL 1
// Core Constants. DO NOT CHANGE
`define IOB_UART_VERSION 16'h0081
