// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_REVERSE_DATA_W 21
// Core Constants. DO NOT CHANGE
`define IOB_REVERSE_VERSION 16'h0081
