// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_XILINX_CLOCK_WIZARD_OUTPUT_PER 1
`define IOB_XILINX_CLOCK_WIZARD_INPUT_PER 1
// Core Constants. DO NOT CHANGE
`define IOB_XILINX_CLOCK_WIZARD_VERSION 16'h0081
