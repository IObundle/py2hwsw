// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_uart_csrs_conf.vh"
`define IOB_CSRS_ADDR_W `IOB_UART_CSRS_ADDR_W
