// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_BOOTROM_AXI_ID_W 1
`define IOB_BOOTROM_AXI_LEN_W 8
// Core Constants. DO NOT CHANGE
`define IOB_BOOTROM_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_BOOTROM_DATA_W 32
`define IOB_BOOTROM_ADDR_W 10
