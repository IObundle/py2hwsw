// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AND_W 21
// Core Constants. DO NOT CHANGE
`define IOB_AND_VERSION 16'h0081
