// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AOI_W 1
// Core Constants. DO NOT CHANGE
`define IOB_AOI_VERSION 16'h0081
