// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXI2IOB_ADDR_WIDTH 32
`define IOB_AXI2IOB_DATA_WIDTH 32
`define IOB_AXI2IOB_STRB_WIDTH (DATA_WIDTH / 8)
`define IOB_AXI2IOB_AXI_ID_WIDTH 8
// Core Constants. DO NOT CHANGE
`define IOB_AXI2IOB_VERSION 16'h0081
