// SPDX-FileCopyrightText: 2024 IObundle
//
// SPDX-License-Identifier: MIT

`define BAUD 115200
`define FREQ 100000000
`define XILINX 1
