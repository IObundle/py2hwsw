// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_UART_TESTER_PBUS_SPLIT_VERSION 16'h0081
