// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_RESET_SYNC_VERSION 16'h0081
