// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_AXI_ID_W 1
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_AXI_LEN_W 4
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_AXI_ADDR_W 28
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_AXI_DATA_W 32
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_BAUD 115200
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_FREQ 50000000
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_MEM_NO_READ_ON_WRITE 1
`define IOB_UART_TESTER_IOB_CYCLONEV_GT_DK_INTEL 1
