// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_RAM_T2P_BE_HEXFILE "none"
`define IOB_RAM_T2P_BE_ADDR_W 1
`define IOB_RAM_T2P_BE_DATA_W 1
// Core Constants. DO NOT CHANGE
`define IOB_RAM_T2P_BE_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_RAM_T2P_BE_COL_W 8
`define IOB_RAM_T2P_BE_NUM_COL DATA_W / COL_W
