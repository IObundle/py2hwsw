// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UNIVERSAL_CONVERTER_AXI_IOB_ADDR_W 1
`define IOB_UNIVERSAL_CONVERTER_AXI_IOB_DATA_W 32
`define IOB_UNIVERSAL_CONVERTER_AXI_IOB_AXI_ID_W 1
`define IOB_UNIVERSAL_CONVERTER_AXI_IOB_AXI_LEN_W 8
// Core Constants. DO NOT CHANGE
`define IOB_UNIVERSAL_CONVERTER_AXI_IOB_VERSION 16'h0081
