// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_IOB2AXIL_AXIL_ADDR_W 21
`define IOB_IOB2AXIL_AXIL_DATA_W 21
`define IOB_IOB2AXIL_ADDR_W AXIL_ADDR_W
`define IOB_IOB2AXIL_DATA_W AXIL_DATA_W
// Core Constants. DO NOT CHANGE
`define IOB_IOB2AXIL_VERSION 16'h0081
