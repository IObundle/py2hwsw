// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UNIVERSAL_CONVERTER_IOB_IOB_ADDR_W 1
`define IOB_UNIVERSAL_CONVERTER_IOB_IOB_DATA_W 32
// Core Constants. DO NOT CHANGE
`define IOB_UNIVERSAL_CONVERTER_IOB_IOB_VERSION 16'h0081
