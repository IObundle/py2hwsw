// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_SYNC_DATA_W 21
`define IOB_SYNC_RST_VAL {DATA_W{1'b0}}
// Core Constants. DO NOT CHANGE
`define IOB_SYNC_VERSION 16'h0081
