//These macros may be dependent on instance parameters
//address macros
//addresses
`define IOB_UART_CSRS_SOFTRESET_ADDR 0
`define IOB_UART_CSRS_SOFTRESET_W 1

`define IOB_UART_CSRS_DIV_ADDR 2
`define IOB_UART_CSRS_DIV_W 16

`define IOB_UART_CSRS_TXDATA_ADDR 4
`define IOB_UART_CSRS_TXDATA_W 8

`define IOB_UART_CSRS_TXEN_ADDR 5
`define IOB_UART_CSRS_TXEN_W 1

`define IOB_UART_CSRS_RXEN_ADDR 6
`define IOB_UART_CSRS_RXEN_W 1

`define IOB_UART_CSRS_TXREADY_ADDR 0
`define IOB_UART_CSRS_TXREADY_W 1

`define IOB_UART_CSRS_RXREADY_ADDR 1
`define IOB_UART_CSRS_RXREADY_W 1

`define IOB_UART_CSRS_RXDATA_ADDR 4
`define IOB_UART_CSRS_RXDATA_W 8

`define IOB_UART_CSRS_VERSION_ADDR 6
`define IOB_UART_CSRS_VERSION_W 16

