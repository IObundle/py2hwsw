// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_REG_CARE_DATA_W 1
`define IOB_REG_CARE_RST_VAL {DATA_W{1'b0}}
// Core Constants. DO NOT CHANGE
`define IOB_REG_CARE_VERSION 16'h0001
