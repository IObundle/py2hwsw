// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_macc_csrs_conf.vh"
`define IOB_CSRS_ADDR_W `IOB_MACC_CSRS_ADDR_W
