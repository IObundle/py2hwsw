// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_TIMER_DATA_W 32
// Core Constants. DO NOT CHANGE
`define IOB_TIMER_VERSION 16'h0081
