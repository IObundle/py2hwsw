// SPDX-FileCopyrightText: 2024 IObundle
//
// SPDX-License-Identifier: MIT

`define BAUD 115200
`define FREQ 50000000
`define INTEL 1
