// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`define IOB_CSRS_ADDR_W axistream_in_csrs_w + axistream_out_csrs_w
